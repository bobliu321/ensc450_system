##
## LEF for PtnCells ;
## created by Innovus v18.10-p002_1 on Tue Apr 20 11:46:48 2021
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ensc450
  CLASS BLOCK ;
  SIZE 375.060000 BY 375.060000 ;
  FOREIGN ensc450 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 156.050000 374.990000 156.120000 375.060000 ;
    END
  END clk
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 155.100000 374.990000 155.170000 375.060000 ;
    END
  END resetn
  PIN EXT_NREADY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 210.035000 375.060000 210.105000 ;
    END
  END EXT_NREADY
  PIN EXT_BUSY
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 219.700000 374.990000 219.770000 375.060000 ;
    END
  END EXT_BUSY
  PIN EXT_MR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 187.400000 374.990000 187.470000 375.060000 ;
    END
  END EXT_MR
  PIN EXT_MW
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 188.350000 374.990000 188.420000 375.060000 ;
    END
  END EXT_MW
  PIN EXT_ADDRBUS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 186.450000 374.990000 186.520000 375.060000 ;
    END
  END EXT_ADDRBUS[31]
  PIN EXT_ADDRBUS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 185.500000 374.990000 185.570000 375.060000 ;
    END
  END EXT_ADDRBUS[30]
  PIN EXT_ADDRBUS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 184.550000 374.990000 184.620000 375.060000 ;
    END
  END EXT_ADDRBUS[29]
  PIN EXT_ADDRBUS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 183.600000 374.990000 183.670000 375.060000 ;
    END
  END EXT_ADDRBUS[28]
  PIN EXT_ADDRBUS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 182.650000 374.990000 182.720000 375.060000 ;
    END
  END EXT_ADDRBUS[27]
  PIN EXT_ADDRBUS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 181.700000 374.990000 181.770000 375.060000 ;
    END
  END EXT_ADDRBUS[26]
  PIN EXT_ADDRBUS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 180.750000 374.990000 180.820000 375.060000 ;
    END
  END EXT_ADDRBUS[25]
  PIN EXT_ADDRBUS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 179.800000 374.990000 179.870000 375.060000 ;
    END
  END EXT_ADDRBUS[24]
  PIN EXT_ADDRBUS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 178.850000 374.990000 178.920000 375.060000 ;
    END
  END EXT_ADDRBUS[23]
  PIN EXT_ADDRBUS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 177.900000 374.990000 177.970000 375.060000 ;
    END
  END EXT_ADDRBUS[22]
  PIN EXT_ADDRBUS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 176.950000 374.990000 177.020000 375.060000 ;
    END
  END EXT_ADDRBUS[21]
  PIN EXT_ADDRBUS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 176.000000 374.990000 176.070000 375.060000 ;
    END
  END EXT_ADDRBUS[20]
  PIN EXT_ADDRBUS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 175.050000 374.990000 175.120000 375.060000 ;
    END
  END EXT_ADDRBUS[19]
  PIN EXT_ADDRBUS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 174.100000 374.990000 174.170000 375.060000 ;
    END
  END EXT_ADDRBUS[18]
  PIN EXT_ADDRBUS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 173.150000 374.990000 173.220000 375.060000 ;
    END
  END EXT_ADDRBUS[17]
  PIN EXT_ADDRBUS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 172.200000 374.990000 172.270000 375.060000 ;
    END
  END EXT_ADDRBUS[16]
  PIN EXT_ADDRBUS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 171.250000 374.990000 171.320000 375.060000 ;
    END
  END EXT_ADDRBUS[15]
  PIN EXT_ADDRBUS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 170.300000 374.990000 170.370000 375.060000 ;
    END
  END EXT_ADDRBUS[14]
  PIN EXT_ADDRBUS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 169.350000 374.990000 169.420000 375.060000 ;
    END
  END EXT_ADDRBUS[13]
  PIN EXT_ADDRBUS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 168.400000 374.990000 168.470000 375.060000 ;
    END
  END EXT_ADDRBUS[12]
  PIN EXT_ADDRBUS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 167.450000 374.990000 167.520000 375.060000 ;
    END
  END EXT_ADDRBUS[11]
  PIN EXT_ADDRBUS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 166.500000 374.990000 166.570000 375.060000 ;
    END
  END EXT_ADDRBUS[10]
  PIN EXT_ADDRBUS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 165.550000 374.990000 165.620000 375.060000 ;
    END
  END EXT_ADDRBUS[9]
  PIN EXT_ADDRBUS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 164.600000 374.990000 164.670000 375.060000 ;
    END
  END EXT_ADDRBUS[8]
  PIN EXT_ADDRBUS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 163.650000 374.990000 163.720000 375.060000 ;
    END
  END EXT_ADDRBUS[7]
  PIN EXT_ADDRBUS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 162.700000 374.990000 162.770000 375.060000 ;
    END
  END EXT_ADDRBUS[6]
  PIN EXT_ADDRBUS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 161.750000 374.990000 161.820000 375.060000 ;
    END
  END EXT_ADDRBUS[5]
  PIN EXT_ADDRBUS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 160.800000 374.990000 160.870000 375.060000 ;
    END
  END EXT_ADDRBUS[4]
  PIN EXT_ADDRBUS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 159.850000 374.990000 159.920000 375.060000 ;
    END
  END EXT_ADDRBUS[3]
  PIN EXT_ADDRBUS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 158.900000 374.990000 158.970000 375.060000 ;
    END
  END EXT_ADDRBUS[2]
  PIN EXT_ADDRBUS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 157.950000 374.990000 158.020000 375.060000 ;
    END
  END EXT_ADDRBUS[1]
  PIN EXT_ADDRBUS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 157.000000 374.990000 157.070000 375.060000 ;
    END
  END EXT_ADDRBUS[0]
  PIN EXT_RDATABUS[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 165.235000 375.060000 165.305000 ;
    END
  END EXT_RDATABUS[31]
  PIN EXT_RDATABUS[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 166.635000 375.060000 166.705000 ;
    END
  END EXT_RDATABUS[30]
  PIN EXT_RDATABUS[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 168.035000 375.060000 168.105000 ;
    END
  END EXT_RDATABUS[29]
  PIN EXT_RDATABUS[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 169.435000 375.060000 169.505000 ;
    END
  END EXT_RDATABUS[28]
  PIN EXT_RDATABUS[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 170.835000 375.060000 170.905000 ;
    END
  END EXT_RDATABUS[27]
  PIN EXT_RDATABUS[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 172.235000 375.060000 172.305000 ;
    END
  END EXT_RDATABUS[26]
  PIN EXT_RDATABUS[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 173.635000 375.060000 173.705000 ;
    END
  END EXT_RDATABUS[25]
  PIN EXT_RDATABUS[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 175.035000 375.060000 175.105000 ;
    END
  END EXT_RDATABUS[24]
  PIN EXT_RDATABUS[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 176.435000 375.060000 176.505000 ;
    END
  END EXT_RDATABUS[23]
  PIN EXT_RDATABUS[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 177.835000 375.060000 177.905000 ;
    END
  END EXT_RDATABUS[22]
  PIN EXT_RDATABUS[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 179.235000 375.060000 179.305000 ;
    END
  END EXT_RDATABUS[21]
  PIN EXT_RDATABUS[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 180.635000 375.060000 180.705000 ;
    END
  END EXT_RDATABUS[20]
  PIN EXT_RDATABUS[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 182.035000 375.060000 182.105000 ;
    END
  END EXT_RDATABUS[19]
  PIN EXT_RDATABUS[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 183.435000 375.060000 183.505000 ;
    END
  END EXT_RDATABUS[18]
  PIN EXT_RDATABUS[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 184.835000 375.060000 184.905000 ;
    END
  END EXT_RDATABUS[17]
  PIN EXT_RDATABUS[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 186.235000 375.060000 186.305000 ;
    END
  END EXT_RDATABUS[16]
  PIN EXT_RDATABUS[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 187.635000 375.060000 187.705000 ;
    END
  END EXT_RDATABUS[15]
  PIN EXT_RDATABUS[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 189.035000 375.060000 189.105000 ;
    END
  END EXT_RDATABUS[14]
  PIN EXT_RDATABUS[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 190.435000 375.060000 190.505000 ;
    END
  END EXT_RDATABUS[13]
  PIN EXT_RDATABUS[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 191.835000 375.060000 191.905000 ;
    END
  END EXT_RDATABUS[12]
  PIN EXT_RDATABUS[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 193.235000 375.060000 193.305000 ;
    END
  END EXT_RDATABUS[11]
  PIN EXT_RDATABUS[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 194.635000 375.060000 194.705000 ;
    END
  END EXT_RDATABUS[10]
  PIN EXT_RDATABUS[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 196.035000 375.060000 196.105000 ;
    END
  END EXT_RDATABUS[9]
  PIN EXT_RDATABUS[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 197.435000 375.060000 197.505000 ;
    END
  END EXT_RDATABUS[8]
  PIN EXT_RDATABUS[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 198.835000 375.060000 198.905000 ;
    END
  END EXT_RDATABUS[7]
  PIN EXT_RDATABUS[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 200.235000 375.060000 200.305000 ;
    END
  END EXT_RDATABUS[6]
  PIN EXT_RDATABUS[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 201.635000 375.060000 201.705000 ;
    END
  END EXT_RDATABUS[5]
  PIN EXT_RDATABUS[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 203.035000 375.060000 203.105000 ;
    END
  END EXT_RDATABUS[4]
  PIN EXT_RDATABUS[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 204.435000 375.060000 204.505000 ;
    END
  END EXT_RDATABUS[3]
  PIN EXT_RDATABUS[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 205.835000 375.060000 205.905000 ;
    END
  END EXT_RDATABUS[2]
  PIN EXT_RDATABUS[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 207.235000 375.060000 207.305000 ;
    END
  END EXT_RDATABUS[1]
  PIN EXT_RDATABUS[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 374.990000 208.635000 375.060000 208.705000 ;
    END
  END EXT_RDATABUS[0]
  PIN EXT_WDATABUS[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 218.750000 374.990000 218.820000 375.060000 ;
    END
  END EXT_WDATABUS[31]
  PIN EXT_WDATABUS[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 217.800000 374.990000 217.870000 375.060000 ;
    END
  END EXT_WDATABUS[30]
  PIN EXT_WDATABUS[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 216.850000 374.990000 216.920000 375.060000 ;
    END
  END EXT_WDATABUS[29]
  PIN EXT_WDATABUS[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 215.900000 374.990000 215.970000 375.060000 ;
    END
  END EXT_WDATABUS[28]
  PIN EXT_WDATABUS[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 214.950000 374.990000 215.020000 375.060000 ;
    END
  END EXT_WDATABUS[27]
  PIN EXT_WDATABUS[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 214.000000 374.990000 214.070000 375.060000 ;
    END
  END EXT_WDATABUS[26]
  PIN EXT_WDATABUS[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 213.050000 374.990000 213.120000 375.060000 ;
    END
  END EXT_WDATABUS[25]
  PIN EXT_WDATABUS[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 212.100000 374.990000 212.170000 375.060000 ;
    END
  END EXT_WDATABUS[24]
  PIN EXT_WDATABUS[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 211.150000 374.990000 211.220000 375.060000 ;
    END
  END EXT_WDATABUS[23]
  PIN EXT_WDATABUS[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 210.200000 374.990000 210.270000 375.060000 ;
    END
  END EXT_WDATABUS[22]
  PIN EXT_WDATABUS[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 209.250000 374.990000 209.320000 375.060000 ;
    END
  END EXT_WDATABUS[21]
  PIN EXT_WDATABUS[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 208.300000 374.990000 208.370000 375.060000 ;
    END
  END EXT_WDATABUS[20]
  PIN EXT_WDATABUS[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 207.350000 374.990000 207.420000 375.060000 ;
    END
  END EXT_WDATABUS[19]
  PIN EXT_WDATABUS[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 206.400000 374.990000 206.470000 375.060000 ;
    END
  END EXT_WDATABUS[18]
  PIN EXT_WDATABUS[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 205.450000 374.990000 205.520000 375.060000 ;
    END
  END EXT_WDATABUS[17]
  PIN EXT_WDATABUS[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 204.500000 374.990000 204.570000 375.060000 ;
    END
  END EXT_WDATABUS[16]
  PIN EXT_WDATABUS[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 203.550000 374.990000 203.620000 375.060000 ;
    END
  END EXT_WDATABUS[15]
  PIN EXT_WDATABUS[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 202.600000 374.990000 202.670000 375.060000 ;
    END
  END EXT_WDATABUS[14]
  PIN EXT_WDATABUS[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 201.650000 374.990000 201.720000 375.060000 ;
    END
  END EXT_WDATABUS[13]
  PIN EXT_WDATABUS[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 200.700000 374.990000 200.770000 375.060000 ;
    END
  END EXT_WDATABUS[12]
  PIN EXT_WDATABUS[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 199.750000 374.990000 199.820000 375.060000 ;
    END
  END EXT_WDATABUS[11]
  PIN EXT_WDATABUS[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 198.800000 374.990000 198.870000 375.060000 ;
    END
  END EXT_WDATABUS[10]
  PIN EXT_WDATABUS[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 197.850000 374.990000 197.920000 375.060000 ;
    END
  END EXT_WDATABUS[9]
  PIN EXT_WDATABUS[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 196.900000 374.990000 196.970000 375.060000 ;
    END
  END EXT_WDATABUS[8]
  PIN EXT_WDATABUS[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 195.950000 374.990000 196.020000 375.060000 ;
    END
  END EXT_WDATABUS[7]
  PIN EXT_WDATABUS[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 195.000000 374.990000 195.070000 375.060000 ;
    END
  END EXT_WDATABUS[6]
  PIN EXT_WDATABUS[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 194.050000 374.990000 194.120000 375.060000 ;
    END
  END EXT_WDATABUS[5]
  PIN EXT_WDATABUS[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 193.100000 374.990000 193.170000 375.060000 ;
    END
  END EXT_WDATABUS[4]
  PIN EXT_WDATABUS[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 192.150000 374.990000 192.220000 375.060000 ;
    END
  END EXT_WDATABUS[3]
  PIN EXT_WDATABUS[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 191.200000 374.990000 191.270000 375.060000 ;
    END
  END EXT_WDATABUS[2]
  PIN EXT_WDATABUS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 190.250000 374.990000 190.320000 375.060000 ;
    END
  END EXT_WDATABUS[1]
  PIN EXT_WDATABUS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 189.300000 374.990000 189.370000 375.060000 ;
    END
  END EXT_WDATABUS[0]
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 375.060000 375.060000 ;
    LAYER metal2 ;
      RECT 219.840000 374.920000 375.060000 375.060000 ;
      RECT 218.890000 374.920000 219.630000 375.060000 ;
      RECT 217.940000 374.920000 218.680000 375.060000 ;
      RECT 216.990000 374.920000 217.730000 375.060000 ;
      RECT 216.040000 374.920000 216.780000 375.060000 ;
      RECT 215.090000 374.920000 215.830000 375.060000 ;
      RECT 214.140000 374.920000 214.880000 375.060000 ;
      RECT 213.190000 374.920000 213.930000 375.060000 ;
      RECT 212.240000 374.920000 212.980000 375.060000 ;
      RECT 211.290000 374.920000 212.030000 375.060000 ;
      RECT 210.340000 374.920000 211.080000 375.060000 ;
      RECT 209.390000 374.920000 210.130000 375.060000 ;
      RECT 208.440000 374.920000 209.180000 375.060000 ;
      RECT 207.490000 374.920000 208.230000 375.060000 ;
      RECT 206.540000 374.920000 207.280000 375.060000 ;
      RECT 205.590000 374.920000 206.330000 375.060000 ;
      RECT 204.640000 374.920000 205.380000 375.060000 ;
      RECT 203.690000 374.920000 204.430000 375.060000 ;
      RECT 202.740000 374.920000 203.480000 375.060000 ;
      RECT 201.790000 374.920000 202.530000 375.060000 ;
      RECT 200.840000 374.920000 201.580000 375.060000 ;
      RECT 199.890000 374.920000 200.630000 375.060000 ;
      RECT 198.940000 374.920000 199.680000 375.060000 ;
      RECT 197.990000 374.920000 198.730000 375.060000 ;
      RECT 197.040000 374.920000 197.780000 375.060000 ;
      RECT 196.090000 374.920000 196.830000 375.060000 ;
      RECT 195.140000 374.920000 195.880000 375.060000 ;
      RECT 194.190000 374.920000 194.930000 375.060000 ;
      RECT 193.240000 374.920000 193.980000 375.060000 ;
      RECT 192.290000 374.920000 193.030000 375.060000 ;
      RECT 191.340000 374.920000 192.080000 375.060000 ;
      RECT 190.390000 374.920000 191.130000 375.060000 ;
      RECT 189.440000 374.920000 190.180000 375.060000 ;
      RECT 188.490000 374.920000 189.230000 375.060000 ;
      RECT 187.540000 374.920000 188.280000 375.060000 ;
      RECT 186.590000 374.920000 187.330000 375.060000 ;
      RECT 185.640000 374.920000 186.380000 375.060000 ;
      RECT 184.690000 374.920000 185.430000 375.060000 ;
      RECT 183.740000 374.920000 184.480000 375.060000 ;
      RECT 182.790000 374.920000 183.530000 375.060000 ;
      RECT 181.840000 374.920000 182.580000 375.060000 ;
      RECT 180.890000 374.920000 181.630000 375.060000 ;
      RECT 179.940000 374.920000 180.680000 375.060000 ;
      RECT 178.990000 374.920000 179.730000 375.060000 ;
      RECT 178.040000 374.920000 178.780000 375.060000 ;
      RECT 177.090000 374.920000 177.830000 375.060000 ;
      RECT 176.140000 374.920000 176.880000 375.060000 ;
      RECT 175.190000 374.920000 175.930000 375.060000 ;
      RECT 174.240000 374.920000 174.980000 375.060000 ;
      RECT 173.290000 374.920000 174.030000 375.060000 ;
      RECT 172.340000 374.920000 173.080000 375.060000 ;
      RECT 171.390000 374.920000 172.130000 375.060000 ;
      RECT 170.440000 374.920000 171.180000 375.060000 ;
      RECT 169.490000 374.920000 170.230000 375.060000 ;
      RECT 168.540000 374.920000 169.280000 375.060000 ;
      RECT 167.590000 374.920000 168.330000 375.060000 ;
      RECT 166.640000 374.920000 167.380000 375.060000 ;
      RECT 165.690000 374.920000 166.430000 375.060000 ;
      RECT 164.740000 374.920000 165.480000 375.060000 ;
      RECT 163.790000 374.920000 164.530000 375.060000 ;
      RECT 162.840000 374.920000 163.580000 375.060000 ;
      RECT 161.890000 374.920000 162.630000 375.060000 ;
      RECT 160.940000 374.920000 161.680000 375.060000 ;
      RECT 159.990000 374.920000 160.730000 375.060000 ;
      RECT 159.040000 374.920000 159.780000 375.060000 ;
      RECT 158.090000 374.920000 158.830000 375.060000 ;
      RECT 157.140000 374.920000 157.880000 375.060000 ;
      RECT 156.190000 374.920000 156.930000 375.060000 ;
      RECT 155.240000 374.920000 155.980000 375.060000 ;
      RECT 0.000000 374.920000 155.030000 375.060000 ;
      RECT 0.000000 210.175000 375.060000 374.920000 ;
      RECT 0.000000 209.965000 374.920000 210.175000 ;
      RECT 0.000000 208.775000 375.060000 209.965000 ;
      RECT 0.000000 208.565000 374.920000 208.775000 ;
      RECT 0.000000 207.375000 375.060000 208.565000 ;
      RECT 0.000000 207.165000 374.920000 207.375000 ;
      RECT 0.000000 205.975000 375.060000 207.165000 ;
      RECT 0.000000 205.765000 374.920000 205.975000 ;
      RECT 0.000000 204.575000 375.060000 205.765000 ;
      RECT 0.000000 204.365000 374.920000 204.575000 ;
      RECT 0.000000 203.175000 375.060000 204.365000 ;
      RECT 0.000000 202.965000 374.920000 203.175000 ;
      RECT 0.000000 201.775000 375.060000 202.965000 ;
      RECT 0.000000 201.565000 374.920000 201.775000 ;
      RECT 0.000000 200.375000 375.060000 201.565000 ;
      RECT 0.000000 200.165000 374.920000 200.375000 ;
      RECT 0.000000 198.975000 375.060000 200.165000 ;
      RECT 0.000000 198.765000 374.920000 198.975000 ;
      RECT 0.000000 197.575000 375.060000 198.765000 ;
      RECT 0.000000 197.365000 374.920000 197.575000 ;
      RECT 0.000000 196.175000 375.060000 197.365000 ;
      RECT 0.000000 195.965000 374.920000 196.175000 ;
      RECT 0.000000 194.775000 375.060000 195.965000 ;
      RECT 0.000000 194.565000 374.920000 194.775000 ;
      RECT 0.000000 193.375000 375.060000 194.565000 ;
      RECT 0.000000 193.165000 374.920000 193.375000 ;
      RECT 0.000000 191.975000 375.060000 193.165000 ;
      RECT 0.000000 191.765000 374.920000 191.975000 ;
      RECT 0.000000 190.575000 375.060000 191.765000 ;
      RECT 0.000000 190.365000 374.920000 190.575000 ;
      RECT 0.000000 189.175000 375.060000 190.365000 ;
      RECT 0.000000 188.965000 374.920000 189.175000 ;
      RECT 0.000000 187.775000 375.060000 188.965000 ;
      RECT 0.000000 187.565000 374.920000 187.775000 ;
      RECT 0.000000 186.375000 375.060000 187.565000 ;
      RECT 0.000000 186.165000 374.920000 186.375000 ;
      RECT 0.000000 184.975000 375.060000 186.165000 ;
      RECT 0.000000 184.765000 374.920000 184.975000 ;
      RECT 0.000000 183.575000 375.060000 184.765000 ;
      RECT 0.000000 183.365000 374.920000 183.575000 ;
      RECT 0.000000 182.175000 375.060000 183.365000 ;
      RECT 0.000000 181.965000 374.920000 182.175000 ;
      RECT 0.000000 180.775000 375.060000 181.965000 ;
      RECT 0.000000 180.565000 374.920000 180.775000 ;
      RECT 0.000000 179.375000 375.060000 180.565000 ;
      RECT 0.000000 179.165000 374.920000 179.375000 ;
      RECT 0.000000 177.975000 375.060000 179.165000 ;
      RECT 0.000000 177.765000 374.920000 177.975000 ;
      RECT 0.000000 176.575000 375.060000 177.765000 ;
      RECT 0.000000 176.365000 374.920000 176.575000 ;
      RECT 0.000000 175.175000 375.060000 176.365000 ;
      RECT 0.000000 174.965000 374.920000 175.175000 ;
      RECT 0.000000 173.775000 375.060000 174.965000 ;
      RECT 0.000000 173.565000 374.920000 173.775000 ;
      RECT 0.000000 172.375000 375.060000 173.565000 ;
      RECT 0.000000 172.165000 374.920000 172.375000 ;
      RECT 0.000000 170.975000 375.060000 172.165000 ;
      RECT 0.000000 170.765000 374.920000 170.975000 ;
      RECT 0.000000 169.575000 375.060000 170.765000 ;
      RECT 0.000000 169.365000 374.920000 169.575000 ;
      RECT 0.000000 168.175000 375.060000 169.365000 ;
      RECT 0.000000 167.965000 374.920000 168.175000 ;
      RECT 0.000000 166.775000 375.060000 167.965000 ;
      RECT 0.000000 166.565000 374.920000 166.775000 ;
      RECT 0.000000 165.375000 375.060000 166.565000 ;
      RECT 0.000000 165.165000 374.920000 165.375000 ;
      RECT 0.000000 0.000000 375.060000 165.165000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 375.060000 375.060000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 375.060000 375.060000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 375.060000 375.060000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 375.060000 375.060000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 375.060000 375.060000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 375.060000 375.060000 ;
    LAYER metal9 ;
      RECT 0.000000 0.000000 375.060000 375.060000 ;
    LAYER metal10 ;
      RECT 0.000000 0.000000 375.060000 375.060000 ;
  END
END ensc450

END LIBRARY
