/local-scratch/localhome/escmc27/ensc450/Project/ensc450_system/syn_045/lib/aesbuffer.lef