##
## LEF for PtnCells ;
## created by Encounter v09.10-p004_1 on Tue Apr  1 17:54:40 2014
##

VERSION 5.5 ;

NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MACRO SRAM
  CLASS BLOCK ;
  SIZE 122.0000 BY 122.0000 ;
  FOREIGN SRAM 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 9.5600 121.9300 9.6300 122.0000 ;
    END
  END clk
  PIN rdn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 10.8900 121.9300 10.9600 122.0000 ;
    END
  END rdn
  PIN wrn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 12.2200 121.9300 12.2900 122.0000 ;
    END
  END wrn
  PIN address[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 26.8500 121.9300 26.9200 122.0000 ;
    END
  END address[10]
  PIN address[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 25.5200 121.9300 25.5900 122.0000 ;
    END
  END address[9]
  PIN address[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 24.1900 121.9300 24.2600 122.0000 ;
    END
  END address[8]
  PIN address[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 22.8600 121.9300 22.9300 122.0000 ;
    END
  END address[7]
  PIN address[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 21.5300 121.9300 21.6000 122.0000 ;
    END
  END address[6]
  PIN address[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 20.2000 121.9300 20.2700 122.0000 ;
    END
  END address[5]
  PIN address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 18.8700 121.9300 18.9400 122.0000 ;
    END
  END address[4]
  PIN address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 17.5400 121.9300 17.6100 122.0000 ;
    END
  END address[3]
  PIN address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 16.2100 121.9300 16.2800 122.0000 ;
    END
  END address[2]
  PIN address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 14.8800 121.9300 14.9500 122.0000 ;
    END
  END address[1]
  PIN address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 13.5500 121.9300 13.6200 122.0000 ;
    END
  END address[0]
  PIN bit_wen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 69.4100 121.9300 69.4800 122.0000 ;
    END
  END bit_wen[31]
  PIN bit_wen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 68.0800 121.9300 68.1500 122.0000 ;
    END
  END bit_wen[30]
  PIN bit_wen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 66.7500 121.9300 66.8200 122.0000 ;
    END
  END bit_wen[29]
  PIN bit_wen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 65.4200 121.9300 65.4900 122.0000 ;
    END
  END bit_wen[28]
  PIN bit_wen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.0900 121.9300 64.1600 122.0000 ;
    END
  END bit_wen[27]
  PIN bit_wen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 62.7600 121.9300 62.8300 122.0000 ;
    END
  END bit_wen[26]
  PIN bit_wen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 61.4300 121.9300 61.5000 122.0000 ;
    END
  END bit_wen[25]
  PIN bit_wen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 60.1000 121.9300 60.1700 122.0000 ;
    END
  END bit_wen[24]
  PIN bit_wen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.7700 121.9300 58.8400 122.0000 ;
    END
  END bit_wen[23]
  PIN bit_wen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 57.4400 121.9300 57.5100 122.0000 ;
    END
  END bit_wen[22]
  PIN bit_wen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 56.1100 121.9300 56.1800 122.0000 ;
    END
  END bit_wen[21]
  PIN bit_wen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 54.7800 121.9300 54.8500 122.0000 ;
    END
  END bit_wen[20]
  PIN bit_wen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 53.4500 121.9300 53.5200 122.0000 ;
    END
  END bit_wen[19]
  PIN bit_wen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.1200 121.9300 52.1900 122.0000 ;
    END
  END bit_wen[18]
  PIN bit_wen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.7900 121.9300 50.8600 122.0000 ;
    END
  END bit_wen[17]
  PIN bit_wen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 49.4600 121.9300 49.5300 122.0000 ;
    END
  END bit_wen[16]
  PIN bit_wen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.1300 121.9300 48.2000 122.0000 ;
    END
  END bit_wen[15]
  PIN bit_wen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 46.8000 121.9300 46.8700 122.0000 ;
    END
  END bit_wen[14]
  PIN bit_wen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 45.4700 121.9300 45.5400 122.0000 ;
    END
  END bit_wen[13]
  PIN bit_wen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 44.1400 121.9300 44.2100 122.0000 ;
    END
  END bit_wen[12]
  PIN bit_wen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 42.8100 121.9300 42.8800 122.0000 ;
    END
  END bit_wen[11]
  PIN bit_wen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 41.4800 121.9300 41.5500 122.0000 ;
    END
  END bit_wen[10]
  PIN bit_wen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 40.1500 121.9300 40.2200 122.0000 ;
    END
  END bit_wen[9]
  PIN bit_wen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 38.8200 121.9300 38.8900 122.0000 ;
    END
  END bit_wen[8]
  PIN bit_wen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 37.4900 121.9300 37.5600 122.0000 ;
    END
  END bit_wen[7]
  PIN bit_wen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 36.1600 121.9300 36.2300 122.0000 ;
    END
  END bit_wen[6]
  PIN bit_wen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 34.8300 121.9300 34.9000 122.0000 ;
    END
  END bit_wen[5]
  PIN bit_wen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.5000 121.9300 33.5700 122.0000 ;
    END
  END bit_wen[4]
  PIN bit_wen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 32.1700 121.9300 32.2400 122.0000 ;
    END
  END bit_wen[3]
  PIN bit_wen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 30.8400 121.9300 30.9100 122.0000 ;
    END
  END bit_wen[2]
  PIN bit_wen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 29.5100 121.9300 29.5800 122.0000 ;
    END
  END bit_wen[1]
  PIN bit_wen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 28.1800 121.9300 28.2500 122.0000 ;
    END
  END bit_wen[0]
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 111.9700 121.9300 112.0400 122.0000 ;
    END
  END data_in[31]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 110.6400 121.9300 110.7100 122.0000 ;
    END
  END data_in[30]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 109.3100 121.9300 109.3800 122.0000 ;
    END
  END data_in[29]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 107.9800 121.9300 108.0500 122.0000 ;
    END
  END data_in[28]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 106.6500 121.9300 106.7200 122.0000 ;
    END
  END data_in[27]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 105.3200 121.9300 105.3900 122.0000 ;
    END
  END data_in[26]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 103.9900 121.9300 104.0600 122.0000 ;
    END
  END data_in[25]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 102.6600 121.9300 102.7300 122.0000 ;
    END
  END data_in[24]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 101.3300 121.9300 101.4000 122.0000 ;
    END
  END data_in[23]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 100.0000 121.9300 100.0700 122.0000 ;
    END
  END data_in[22]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 98.6700 121.9300 98.7400 122.0000 ;
    END
  END data_in[21]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 97.3400 121.9300 97.4100 122.0000 ;
    END
  END data_in[20]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 96.0100 121.9300 96.0800 122.0000 ;
    END
  END data_in[19]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 94.6800 121.9300 94.7500 122.0000 ;
    END
  END data_in[18]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 93.3500 121.9300 93.4200 122.0000 ;
    END
  END data_in[17]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 92.0200 121.9300 92.0900 122.0000 ;
    END
  END data_in[16]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 90.6900 121.9300 90.7600 122.0000 ;
    END
  END data_in[15]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 89.3600 121.9300 89.4300 122.0000 ;
    END
  END data_in[14]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 88.0300 121.9300 88.1000 122.0000 ;
    END
  END data_in[13]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 86.7000 121.9300 86.7700 122.0000 ;
    END
  END data_in[12]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 85.3700 121.9300 85.4400 122.0000 ;
    END
  END data_in[11]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 84.0400 121.9300 84.1100 122.0000 ;
    END
  END data_in[10]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 82.7100 121.9300 82.7800 122.0000 ;
    END
  END data_in[9]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 81.3800 121.9300 81.4500 122.0000 ;
    END
  END data_in[8]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 80.0500 121.9300 80.1200 122.0000 ;
    END
  END data_in[7]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 78.7200 121.9300 78.7900 122.0000 ;
    END
  END data_in[6]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 77.3900 121.9300 77.4600 122.0000 ;
    END
  END data_in[5]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 76.0600 121.9300 76.1300 122.0000 ;
    END
  END data_in[4]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 74.7300 121.9300 74.8000 122.0000 ;
    END
  END data_in[3]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 73.4000 121.9300 73.4700 122.0000 ;
    END
  END data_in[2]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 72.0700 121.9300 72.1400 122.0000 ;
    END
  END data_in[1]
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 70.7400 121.9300 70.8100 122.0000 ;
    END
  END data_in[0]
  PIN data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 93.2750 122.0000 93.3450 ;
    END
  END data_out[31]
  PIN data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 91.1750 122.0000 91.2450 ;
    END
  END data_out[30]
  PIN data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 89.0750 122.0000 89.1450 ;
    END
  END data_out[29]
  PIN data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 86.9750 122.0000 87.0450 ;
    END
  END data_out[28]
  PIN data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 84.8750 122.0000 84.9450 ;
    END
  END data_out[27]
  PIN data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 82.7750 122.0000 82.8450 ;
    END
  END data_out[26]
  PIN data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 80.6750 122.0000 80.7450 ;
    END
  END data_out[25]
  PIN data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 78.5750 122.0000 78.6450 ;
    END
  END data_out[24]
  PIN data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 76.4750 122.0000 76.5450 ;
    END
  END data_out[23]
  PIN data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 74.3750 122.0000 74.4450 ;
    END
  END data_out[22]
  PIN data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 72.2750 122.0000 72.3450 ;
    END
  END data_out[21]
  PIN data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 70.1750 122.0000 70.2450 ;
    END
  END data_out[20]
  PIN data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 68.0750 122.0000 68.1450 ;
    END
  END data_out[19]
  PIN data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 65.9750 122.0000 66.0450 ;
    END
  END data_out[18]
  PIN data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 63.8750 122.0000 63.9450 ;
    END
  END data_out[17]
  PIN data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 61.7750 122.0000 61.8450 ;
    END
  END data_out[16]
  PIN data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 59.6750 122.0000 59.7450 ;
    END
  END data_out[15]
  PIN data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 57.5750 122.0000 57.6450 ;
    END
  END data_out[14]
  PIN data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 55.4750 122.0000 55.5450 ;
    END
  END data_out[13]
  PIN data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 53.3750 122.0000 53.4450 ;
    END
  END data_out[12]
  PIN data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 51.2750 122.0000 51.3450 ;
    END
  END data_out[11]
  PIN data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 49.1750 122.0000 49.2450 ;
    END
  END data_out[10]
  PIN data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 47.0750 122.0000 47.1450 ;
    END
  END data_out[9]
  PIN data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 44.9750 122.0000 45.0450 ;
    END
  END data_out[8]
  PIN data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 42.8750 122.0000 42.9450 ;
    END
  END data_out[7]
  PIN data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 40.7750 122.0000 40.8450 ;
    END
  END data_out[6]
  PIN data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 38.6750 122.0000 38.7450 ;
    END
  END data_out[5]
  PIN data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 36.5750 122.0000 36.6450 ;
    END
  END data_out[4]
  PIN data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 34.4750 122.0000 34.5450 ;
    END
  END data_out[3]
  PIN data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 32.3750 122.0000 32.4450 ;
    END
  END data_out[2]
  PIN data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 30.2750 122.0000 30.3450 ;
    END
  END data_out[1]
  PIN data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 121.9300 28.1750 122.0000 28.2450 ;
    END
  END data_out[0]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal10 ;
        RECT 2.3800 0.0000 3.1800 0.8000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 2.3800 121.2000 3.1800 122.0000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 118.9900 0.0000 119.7900 0.8000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 118.9900 121.2000 119.7900 122.0000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal10 ;
        RECT 0.7800 0.0000 1.5800 0.8000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 0.7800 121.2000 1.5800 122.0000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 120.5900 0.0000 121.3900 0.8000 ;
    END
    PORT
      LAYER metal10 ;
        RECT 120.5900 121.2000 121.3900 122.0000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.0000 0.0000 122.0000 122.0000 ;
    LAYER metal2 ;
      RECT 112.1100 121.8600 122.0000 122.0000 ;
      RECT 110.7800 121.8600 111.9000 122.0000 ;
      RECT 109.4500 121.8600 110.5700 122.0000 ;
      RECT 108.1200 121.8600 109.2400 122.0000 ;
      RECT 106.7900 121.8600 107.9100 122.0000 ;
      RECT 105.4600 121.8600 106.5800 122.0000 ;
      RECT 104.1300 121.8600 105.2500 122.0000 ;
      RECT 102.8000 121.8600 103.9200 122.0000 ;
      RECT 101.4700 121.8600 102.5900 122.0000 ;
      RECT 100.1400 121.8600 101.2600 122.0000 ;
      RECT 98.8100 121.8600 99.9300 122.0000 ;
      RECT 97.4800 121.8600 98.6000 122.0000 ;
      RECT 96.1500 121.8600 97.2700 122.0000 ;
      RECT 94.8200 121.8600 95.9400 122.0000 ;
      RECT 93.4900 121.8600 94.6100 122.0000 ;
      RECT 92.1600 121.8600 93.2800 122.0000 ;
      RECT 90.8300 121.8600 91.9500 122.0000 ;
      RECT 89.5000 121.8600 90.6200 122.0000 ;
      RECT 88.1700 121.8600 89.2900 122.0000 ;
      RECT 86.8400 121.8600 87.9600 122.0000 ;
      RECT 85.5100 121.8600 86.6300 122.0000 ;
      RECT 84.1800 121.8600 85.3000 122.0000 ;
      RECT 82.8500 121.8600 83.9700 122.0000 ;
      RECT 81.5200 121.8600 82.6400 122.0000 ;
      RECT 80.1900 121.8600 81.3100 122.0000 ;
      RECT 78.8600 121.8600 79.9800 122.0000 ;
      RECT 77.5300 121.8600 78.6500 122.0000 ;
      RECT 76.2000 121.8600 77.3200 122.0000 ;
      RECT 74.8700 121.8600 75.9900 122.0000 ;
      RECT 73.5400 121.8600 74.6600 122.0000 ;
      RECT 72.2100 121.8600 73.3300 122.0000 ;
      RECT 70.8800 121.8600 72.0000 122.0000 ;
      RECT 69.5500 121.8600 70.6700 122.0000 ;
      RECT 68.2200 121.8600 69.3400 122.0000 ;
      RECT 66.8900 121.8600 68.0100 122.0000 ;
      RECT 65.5600 121.8600 66.6800 122.0000 ;
      RECT 64.2300 121.8600 65.3500 122.0000 ;
      RECT 62.9000 121.8600 64.0200 122.0000 ;
      RECT 61.5700 121.8600 62.6900 122.0000 ;
      RECT 60.2400 121.8600 61.3600 122.0000 ;
      RECT 58.9100 121.8600 60.0300 122.0000 ;
      RECT 57.5800 121.8600 58.7000 122.0000 ;
      RECT 56.2500 121.8600 57.3700 122.0000 ;
      RECT 54.9200 121.8600 56.0400 122.0000 ;
      RECT 53.5900 121.8600 54.7100 122.0000 ;
      RECT 52.2600 121.8600 53.3800 122.0000 ;
      RECT 50.9300 121.8600 52.0500 122.0000 ;
      RECT 49.6000 121.8600 50.7200 122.0000 ;
      RECT 48.2700 121.8600 49.3900 122.0000 ;
      RECT 46.9400 121.8600 48.0600 122.0000 ;
      RECT 45.6100 121.8600 46.7300 122.0000 ;
      RECT 44.2800 121.8600 45.4000 122.0000 ;
      RECT 42.9500 121.8600 44.0700 122.0000 ;
      RECT 41.6200 121.8600 42.7400 122.0000 ;
      RECT 40.2900 121.8600 41.4100 122.0000 ;
      RECT 38.9600 121.8600 40.0800 122.0000 ;
      RECT 37.6300 121.8600 38.7500 122.0000 ;
      RECT 36.3000 121.8600 37.4200 122.0000 ;
      RECT 34.9700 121.8600 36.0900 122.0000 ;
      RECT 33.6400 121.8600 34.7600 122.0000 ;
      RECT 32.3100 121.8600 33.4300 122.0000 ;
      RECT 30.9800 121.8600 32.1000 122.0000 ;
      RECT 29.6500 121.8600 30.7700 122.0000 ;
      RECT 28.3200 121.8600 29.4400 122.0000 ;
      RECT 26.9900 121.8600 28.1100 122.0000 ;
      RECT 25.6600 121.8600 26.7800 122.0000 ;
      RECT 24.3300 121.8600 25.4500 122.0000 ;
      RECT 23.0000 121.8600 24.1200 122.0000 ;
      RECT 21.6700 121.8600 22.7900 122.0000 ;
      RECT 20.3400 121.8600 21.4600 122.0000 ;
      RECT 19.0100 121.8600 20.1300 122.0000 ;
      RECT 17.6800 121.8600 18.8000 122.0000 ;
      RECT 16.3500 121.8600 17.4700 122.0000 ;
      RECT 15.0200 121.8600 16.1400 122.0000 ;
      RECT 13.6900 121.8600 14.8100 122.0000 ;
      RECT 12.3600 121.8600 13.4800 122.0000 ;
      RECT 11.0300 121.8600 12.1500 122.0000 ;
      RECT 9.7000 121.8600 10.8200 122.0000 ;
      RECT 0.0000 121.8600 9.4900 122.0000 ;
      RECT 0.0000 93.4150 122.0000 121.8600 ;
      RECT 0.0000 93.2050 121.8600 93.4150 ;
      RECT 0.0000 91.3150 122.0000 93.2050 ;
      RECT 0.0000 91.1050 121.8600 91.3150 ;
      RECT 0.0000 89.2150 122.0000 91.1050 ;
      RECT 0.0000 89.0050 121.8600 89.2150 ;
      RECT 0.0000 87.1150 122.0000 89.0050 ;
      RECT 0.0000 86.9050 121.8600 87.1150 ;
      RECT 0.0000 85.0150 122.0000 86.9050 ;
      RECT 0.0000 84.8050 121.8600 85.0150 ;
      RECT 0.0000 82.9150 122.0000 84.8050 ;
      RECT 0.0000 82.7050 121.8600 82.9150 ;
      RECT 0.0000 80.8150 122.0000 82.7050 ;
      RECT 0.0000 80.6050 121.8600 80.8150 ;
      RECT 0.0000 78.7150 122.0000 80.6050 ;
      RECT 0.0000 78.5050 121.8600 78.7150 ;
      RECT 0.0000 76.6150 122.0000 78.5050 ;
      RECT 0.0000 76.4050 121.8600 76.6150 ;
      RECT 0.0000 74.5150 122.0000 76.4050 ;
      RECT 0.0000 74.3050 121.8600 74.5150 ;
      RECT 0.0000 72.4150 122.0000 74.3050 ;
      RECT 0.0000 72.2050 121.8600 72.4150 ;
      RECT 0.0000 70.3150 122.0000 72.2050 ;
      RECT 0.0000 70.1050 121.8600 70.3150 ;
      RECT 0.0000 68.2150 122.0000 70.1050 ;
      RECT 0.0000 68.0050 121.8600 68.2150 ;
      RECT 0.0000 66.1150 122.0000 68.0050 ;
      RECT 0.0000 65.9050 121.8600 66.1150 ;
      RECT 0.0000 64.0150 122.0000 65.9050 ;
      RECT 0.0000 63.8050 121.8600 64.0150 ;
      RECT 0.0000 61.9150 122.0000 63.8050 ;
      RECT 0.0000 61.7050 121.8600 61.9150 ;
      RECT 0.0000 59.8150 122.0000 61.7050 ;
      RECT 0.0000 59.6050 121.8600 59.8150 ;
      RECT 0.0000 57.7150 122.0000 59.6050 ;
      RECT 0.0000 57.5050 121.8600 57.7150 ;
      RECT 0.0000 55.6150 122.0000 57.5050 ;
      RECT 0.0000 55.4050 121.8600 55.6150 ;
      RECT 0.0000 53.5150 122.0000 55.4050 ;
      RECT 0.0000 53.3050 121.8600 53.5150 ;
      RECT 0.0000 51.4150 122.0000 53.3050 ;
      RECT 0.0000 51.2050 121.8600 51.4150 ;
      RECT 0.0000 49.3150 122.0000 51.2050 ;
      RECT 0.0000 49.1050 121.8600 49.3150 ;
      RECT 0.0000 47.2150 122.0000 49.1050 ;
      RECT 0.0000 47.0050 121.8600 47.2150 ;
      RECT 0.0000 45.1150 122.0000 47.0050 ;
      RECT 0.0000 44.9050 121.8600 45.1150 ;
      RECT 0.0000 43.0150 122.0000 44.9050 ;
      RECT 0.0000 42.8050 121.8600 43.0150 ;
      RECT 0.0000 40.9150 122.0000 42.8050 ;
      RECT 0.0000 40.7050 121.8600 40.9150 ;
      RECT 0.0000 38.8150 122.0000 40.7050 ;
      RECT 0.0000 38.6050 121.8600 38.8150 ;
      RECT 0.0000 36.7150 122.0000 38.6050 ;
      RECT 0.0000 36.5050 121.8600 36.7150 ;
      RECT 0.0000 34.6150 122.0000 36.5050 ;
      RECT 0.0000 34.4050 121.8600 34.6150 ;
      RECT 0.0000 32.5150 122.0000 34.4050 ;
      RECT 0.0000 32.3050 121.8600 32.5150 ;
      RECT 0.0000 30.4150 122.0000 32.3050 ;
      RECT 0.0000 30.2050 121.8600 30.4150 ;
      RECT 0.0000 28.3150 122.0000 30.2050 ;
      RECT 0.0000 28.1050 121.8600 28.3150 ;
      RECT 0.0000 0.0000 122.0000 28.1050 ;
    LAYER metal3 ;
      RECT 0.0000 0.0000 122.0000 122.0000 ;
    LAYER metal4 ;
      RECT 0.0000 0.0000 122.0000 122.0000 ;
  END
END SRAM

END LIBRARY
