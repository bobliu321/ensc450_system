/local-scratch/localhome/escmc27/ensc450/Project/ensc450_system/vhdl/SRAM_Lib/SRAM.lef